magic
tech scmos
timestamp 1591015897
<< error_p >>
rect -14 9 16 11
rect -14 8 15 9
rect -13 7 -9 8
rect -13 6 0 7
rect 9 6 15 7
rect -13 5 -10 6
rect -6 5 -3 6
rect 1 5 4 6
rect 12 5 15 6
rect -13 4 15 5
rect -13 2 -6 4
rect -3 2 -2 4
rect 4 2 5 4
rect 15 2 16 4
rect -14 -1 16 1
rect -17 -9 -7 -7
rect -6 -8 -4 -6
rect -6 -9 3 -8
rect -17 -11 0 -9
rect -17 -13 7 -11
rect -16 -14 -7 -13
rect 12 -14 15 -13
rect -13 -15 15 -14
rect -10 -17 -9 -15
rect 15 -17 16 -15
rect -13 -21 -10 -19
rect -10 -23 -9 -21
<< nwell >>
rect -14 1 16 9
<< polysilicon >>
rect -9 4 -7 9
rect -2 4 0 9
rect 5 4 7 9
rect -9 -15 -7 2
rect -2 -15 0 2
rect 5 -15 7 2
rect -9 -19 -7 -17
rect -2 -19 0 -17
rect 5 -19 7 -17
<< ndiffusion >>
rect -10 -17 -9 -15
rect -7 -17 -2 -15
rect 0 -17 5 -15
rect 7 -17 12 -15
<< pdiffusion >>
rect -10 2 -9 4
rect -7 2 -6 4
rect -3 2 -2 4
rect 0 2 1 4
rect 4 2 5 4
rect 7 2 12 4
<< metal1 >>
rect -14 6 -13 8
rect -10 6 15 8
rect -13 4 -10 6
rect 1 4 4 6
rect -6 -6 -3 2
rect 12 -6 15 2
rect -6 -9 15 -6
rect -17 -10 -7 -9
rect -17 -12 0 -11
rect -17 -14 7 -13
rect 12 -15 15 -9
rect -13 -20 -10 -17
rect -13 -21 15 -20
rect -10 -23 15 -21
<< ntransistor >>
rect -9 -17 -7 -15
rect -2 -17 0 -15
rect 5 -17 7 -15
<< ptransistor >>
rect -9 2 -7 4
rect -2 2 0 4
rect 5 2 7 4
<< ndcontact >>
rect -13 -17 -10 -15
rect 12 -17 15 -15
<< pdcontact >>
rect -13 2 -10 4
rect -6 2 -3 4
rect 1 2 4 4
rect 12 2 15 4
<< psubstratepcontact >>
rect -13 -23 -10 -21
<< nsubstratencontact >>
rect -13 6 -10 8
<< labels >>
rlabel metal1 -5 7 -5 7 5 Vdd!
rlabel metal1 -4 -22 -4 -22 1 Gnd!
rlabel ndiffusion 3 -16 3 -16 1 ntype+
rlabel pdiffusion 9 3 9 3 1 ptype+
rlabel metal1 -17 -10 -17 -10 3 input1+
rlabel metal1 -17 -12 -17 -12 3 input2+
rlabel metal1 -17 -14 -17 -14 3 input3+
<< end >>
